module add1(
	input a,b,c,
	output s,co
);
assign s=(c+a+b);
assign co=(c+a+b);

endmodule